`timescale 1ns / 1ps


module router_top(
    input clk,
    input resetn,
    input packet_valid,
    // Read enables from the external receivers for each output channel
    input read_enb_0,
    input read_enb_1,
    input read_enb_2,
    input [7:0] datain,

    output vldout_0, vldout_1, vldout_2, // Valid signals for each output channel
    output err,      // Parity error flag
    output busy,     // Router busy flag
    output [7:0] data_out_0, data_out_1, data_out_2 // Data outputs for each channel
);


    // Control signals generated by the FSM
    wire detect_add, ld_state, laf_state, lfd_state, full_state, rst_int_reg, write_enb_reg;

    // Status signals generated by the Register module
    wire err, parity_done, low_packet_valid;

    // Data output from the Register module, which feeds into the FIFOs
    wire [7:0] dout;

    // Status signals from the Synchronizer to the FSM
    wire fifo_full;

    // Control signals from the Synchronizer to the FIFOs
    wire [2:0] w_enb;       // 3-bit write enable for the three FIFOs
    wire [2:0] soft_reset;  // 3-bit soft reset for the three FIFOs

    // Status signals from the three FIFOs to the Synchronizer
    wire [2:0] empty;       // 3-bit empty status
    wire [2:0] full;        // 3-bit full status

    // Temporary wire array to hold the data outputs from the three FIFOs
    wire [7:0] data_out_temp[2:0];


    genvar a;
    generate
        for(a=0; a<3; a=a+1) begin: fifo_instance
            // NOTE: The port names below have been updated to match your new router_fifo module.
            router_fifo fifo (
                .clk(clk),
                .resetn(resetn),
                .soft_reset(soft_reset[a]),
                .lfd_state(lfd_state),
                .wr_en(w_enb[a]),           // Changed from .write_enb
                .data_in(dout),             // Changed from .datain
                .rd_en( (a==0) ? read_enb_0 : (a==1) ? read_enb_1 : read_enb_2 ), // Changed from .read_enb
                .full(full[a]),
                .empty(empty[a]),
                .data_out(data_out_temp[a]) // Changed from .dataout
            );
        end
    endgenerate


    router_register r1 (
        .clk(clk),
        .resetn(resetn),
        .packet_valid(packet_valid),
        .datain(datain),
        .fifo_full(fifo_full), // Gets full status from the Synchronizer
        .detect_add(detect_add),
        .ld_state(ld_state),
        .laf_state(laf_state),
        .full_state(full_state),
        .lfd_state(lfd_state),
        .rst_int_reg(rst_int_reg),
        .dout(dout), 
        .err(err),
        .parity_done(parity_done),
        .low_packet_valid(low_packet_valid)
    );

    router_fsm fsm (
        .clk(clk),
        .resetn(resetn),
        .packet_valid(packet_valid),
        .datain(datain[1:0]), // FSM only needs the 2 address bits from datain
        .fifo_full(fifo_full),
        .fifo_empty_0(empty[0]),
        .fifo_empty_1(empty[1]),
        .fifo_empty_2(empty[2]),
        .soft_reset_0(soft_reset[0]),
        .soft_reset_1(soft_reset[1]),
        .soft_reset_2(soft_reset[2]),
        .parity_done(parity_done),
        .low_packet_valid(low_packet_valid),
        .busy(busy),
        .rst_int_reg(rst_int_reg),
        .full_state(full_state),
        .lfd_state(lfd_state),
        .laf_state(laf_state),
        .ld_state(ld_state),
        .detect_add(detect_add),
        .write_enb_reg(write_enb_reg)
    );

    router_synchronizer sync (
        .clk(clk),
        .resetn(resetn),
        .datain(datain[1:0]), // Sync also needs the 2 address bits
        .detect_add(detect_add),
        .write_enb_reg(write_enb_reg),
        .full_0(full[0]), .full_1(full[1]), .full_2(full[2]),
        .empty_0(empty[0]), .empty_1(empty[1]), .empty_2(empty[2]),
        .read_enb_0(read_enb_0), .read_enb_1(read_enb_1), .read_enb_2(read_enb_2),
        .vld_out_0(vldout_0), .vld_out_1(vldout_1), .vld_out_2(vldout_2),
        .soft_reset_0(soft_reset[0]), .soft_reset_1(soft_reset[1]), .soft_reset_2(soft_reset[2]),
        .write_enb(w_enb),
        .fifo_full(fifo_full)
    );


    assign data_out_0 = data_out_temp[0];
    assign data_out_1 = data_out_temp[1];
    assign data_out_2 = data_out_temp[2];

endmodule

